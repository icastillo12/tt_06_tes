VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_inverter
  CLASS BLOCK ;
  FOREIGN tt_um_inverter ;
  ORIGIN -1.000 0.100 ;
  SIZE 157.900 BY 226.470 ;
  OBS
      LAYER nwell ;
        RECT 27.370 10.675 28.410 12.215 ;
      LAYER pwell ;
        RECT 27.420 8.920 28.360 10.240 ;
      LAYER li1 ;
        RECT 27.560 11.755 28.220 12.025 ;
        RECT 27.590 10.855 27.760 11.755 ;
        RECT 27.625 10.305 27.795 10.635 ;
        RECT 28.020 10.585 28.190 11.405 ;
        RECT 28.020 10.415 29.230 10.585 ;
        RECT 27.590 9.330 27.760 10.110 ;
        RECT 28.020 9.690 28.190 10.415 ;
        RECT 27.560 9.060 28.220 9.330 ;
      LAYER mcon ;
        RECT 27.805 11.805 27.975 11.975 ;
        RECT 27.625 10.385 27.795 10.555 ;
        RECT 28.980 10.415 29.150 10.585 ;
        RECT 27.805 9.110 27.975 9.280 ;
      LAYER met1 ;
        RECT 27.190 11.750 28.590 12.120 ;
        RECT 27.595 10.540 27.825 10.615 ;
        RECT 10.305 10.400 27.825 10.540 ;
        RECT 10.305 3.060 10.445 10.400 ;
        RECT 27.595 10.325 27.825 10.400 ;
        RECT 28.885 10.345 32.700 10.650 ;
        RECT 29.265 10.340 32.700 10.345 ;
        RECT 27.275 8.965 28.675 9.335 ;
        RECT 2.095 2.920 10.445 3.060 ;
        RECT 24.090 2.930 24.370 3.215 ;
        RECT 32.390 2.930 32.700 10.340 ;
        RECT 2.095 1.490 2.375 2.920 ;
        RECT 24.090 2.620 32.700 2.930 ;
        RECT 24.090 1.645 24.370 2.620 ;
      LAYER via ;
        RECT 27.280 11.805 27.540 12.065 ;
        RECT 27.600 11.805 27.860 12.065 ;
        RECT 27.920 11.805 28.180 12.065 ;
        RECT 28.240 11.805 28.500 12.065 ;
        RECT 27.365 9.020 27.625 9.280 ;
        RECT 27.685 9.020 27.945 9.280 ;
        RECT 28.005 9.020 28.265 9.280 ;
        RECT 28.325 9.020 28.585 9.280 ;
        RECT 2.105 2.625 2.365 2.885 ;
        RECT 2.105 2.305 2.365 2.565 ;
        RECT 2.105 1.985 2.365 2.245 ;
        RECT 2.105 1.665 2.365 1.925 ;
        RECT 24.100 2.780 24.360 3.040 ;
        RECT 24.100 2.460 24.360 2.720 ;
        RECT 24.100 2.140 24.360 2.400 ;
        RECT 24.100 1.820 24.360 2.080 ;
      LAYER met2 ;
        RECT 27.190 11.750 28.590 12.120 ;
        RECT 27.275 8.965 28.675 9.335 ;
        RECT 2.095 1.490 2.375 3.060 ;
        RECT 24.090 1.645 24.370 3.215 ;
      LAYER via2 ;
        RECT 27.350 11.795 27.630 12.075 ;
        RECT 27.750 11.795 28.030 12.075 ;
        RECT 28.150 11.795 28.430 12.075 ;
        RECT 27.435 9.010 27.715 9.290 ;
        RECT 27.835 9.010 28.115 9.290 ;
        RECT 28.235 9.010 28.515 9.290 ;
        RECT 2.095 2.735 2.375 3.015 ;
        RECT 2.095 2.335 2.375 2.615 ;
        RECT 2.095 1.935 2.375 2.215 ;
        RECT 2.095 1.535 2.375 1.815 ;
        RECT 24.090 2.890 24.370 3.170 ;
        RECT 24.090 2.490 24.370 2.770 ;
        RECT 24.090 2.090 24.370 2.370 ;
        RECT 24.090 1.690 24.370 1.970 ;
      LAYER met3 ;
        RECT 27.130 11.745 28.650 12.125 ;
        RECT 27.215 8.960 28.735 9.340 ;
        RECT 2.070 1.485 2.400 3.065 ;
        RECT 24.065 1.640 24.395 3.220 ;
      LAYER via3 ;
        RECT 27.130 11.775 27.450 12.095 ;
        RECT 27.530 11.775 27.850 12.095 ;
        RECT 27.930 11.775 28.250 12.095 ;
        RECT 28.330 11.775 28.650 12.095 ;
        RECT 27.215 8.990 27.535 9.310 ;
        RECT 27.615 8.990 27.935 9.310 ;
        RECT 28.015 8.990 28.335 9.310 ;
        RECT 28.415 8.990 28.735 9.310 ;
        RECT 2.075 2.715 2.395 3.035 ;
        RECT 2.075 2.315 2.395 2.635 ;
        RECT 2.075 1.915 2.395 2.235 ;
        RECT 2.075 1.515 2.395 1.835 ;
        RECT 24.070 2.870 24.390 3.190 ;
        RECT 24.070 2.470 24.390 2.790 ;
        RECT 24.070 2.070 24.390 2.390 ;
        RECT 24.070 1.670 24.390 1.990 ;
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
        RECT 7.670 224.760 7.970 225.760 ;
        RECT 11.350 224.760 11.650 225.760 ;
        RECT 15.030 224.760 15.330 225.760 ;
        RECT 18.710 224.760 19.010 225.760 ;
        RECT 22.390 224.760 22.690 225.760 ;
        RECT 26.070 224.760 26.370 225.760 ;
        RECT 29.750 224.760 30.050 225.760 ;
        RECT 33.430 224.760 33.730 225.760 ;
        RECT 37.110 224.760 37.410 225.760 ;
        RECT 40.790 224.760 41.090 225.760 ;
        RECT 44.470 224.760 44.770 225.760 ;
        RECT 48.150 224.760 48.450 225.760 ;
        RECT 51.830 224.760 52.130 225.760 ;
        RECT 55.510 224.760 55.810 225.760 ;
        RECT 59.190 224.760 59.490 225.760 ;
        RECT 62.870 224.760 63.170 225.760 ;
        RECT 66.550 224.760 66.850 225.760 ;
        RECT 70.230 224.760 70.530 225.760 ;
        RECT 73.910 224.760 74.210 225.760 ;
        RECT 77.590 224.760 77.890 225.760 ;
        RECT 81.270 224.760 81.570 225.760 ;
        RECT 84.950 224.760 85.250 225.760 ;
        RECT 88.630 224.760 88.930 225.760 ;
        RECT 92.310 224.760 92.610 225.760 ;
        RECT 95.990 224.760 96.290 225.760 ;
        RECT 99.670 224.760 99.970 225.760 ;
        RECT 103.350 224.760 103.650 225.760 ;
        RECT 107.030 224.760 107.330 225.760 ;
        RECT 110.710 224.760 111.010 225.760 ;
        RECT 114.390 224.760 114.690 225.760 ;
        RECT 118.070 224.760 118.370 225.760 ;
        RECT 121.750 224.760 122.050 225.760 ;
        RECT 125.430 224.760 125.730 225.760 ;
        RECT 129.110 224.760 129.410 225.760 ;
        RECT 132.790 224.760 133.090 225.760 ;
        RECT 136.470 224.760 136.770 225.760 ;
        RECT 140.150 224.760 140.450 225.760 ;
        RECT 143.830 224.760 144.130 225.760 ;
        RECT 147.510 224.760 147.810 225.760 ;
        RECT 151.190 224.760 151.490 225.760 ;
        RECT 154.870 224.760 155.170 225.760 ;
        RECT 158.550 224.760 158.850 225.760 ;
        RECT 1.000 12.085 2.500 220.760 ;
        RECT 27.125 12.085 28.655 12.100 ;
        RECT 1.000 11.785 28.655 12.085 ;
        RECT 1.000 5.000 2.500 11.785 ;
        RECT 27.125 11.770 28.655 11.785 ;
        RECT 27.210 9.300 28.740 9.315 ;
        RECT 49.000 9.300 50.500 220.760 ;
        RECT 27.210 9.000 50.500 9.300 ;
        RECT 27.210 8.985 28.740 9.000 ;
        RECT 49.000 5.000 50.500 9.000 ;
        RECT 2.070 1.510 2.400 3.040 ;
        RECT 24.065 1.665 24.395 3.195 ;
        RECT 2.070 1.000 2.370 1.510 ;
        RECT 24.095 1.000 24.395 1.665 ;
        RECT 2.000 0.000 2.600 1.000 ;
        RECT 24.080 0.000 24.680 1.000 ;
        RECT 46.160 0.000 46.760 1.000 ;
        RECT 68.240 0.000 68.840 1.000 ;
        RECT 90.320 0.000 90.920 1.000 ;
        RECT 112.400 0.000 113.000 1.000 ;
        RECT 134.480 0.000 135.080 1.000 ;
        RECT 156.560 0.000 157.160 1.000 ;
  END
END tt_um_inverter
END LIBRARY

